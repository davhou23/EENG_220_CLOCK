module EENG_220_PROJECT();


endmodule 