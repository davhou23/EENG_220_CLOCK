module EENG_220_PROJECT();

    //HI
endmodule 